BZh91AY&SYM[�X _�Py����߰?���P[А"P�sbh0�2d��`�i���!����a2dɑ��4�# C �!
&�o)�~�b d������a2dɑ��4�# C T�&ѦH(m2M2 40L��M���I)t#"^�0% ���jE"��"R�UC��%�M#���0�a�-�۽G��1�ϟ:��pG��	����^���65���ۅ���l<��'"D�"��n}���� <,X'�x�85�a͠>Ql�̤�4gbF|�3G��æe���JU{�{���L�HU7;nM����b�N�>|UW�q�w���+���Fa(�E�®Z�)�pck�0��}�H��]b�c�����A��h�-k��e���\�ƞͱ�m@�.a�A�/�k>4L�vZԟtx�"S�d�������s��a`�E�/5��T0S���1Ѝlw)$��!MX�ѭ�c|Y��y��%��1~]'���Լ�p�?�{</R���bY�%�R_�����������Z�R�З�u|=vٚX٭��&�Y���h���$�I����!)Vu�O:�ji��;Sr�Cv�ަ��#_Z�O	��ꪓ�Ћ't�ƒM�'.�R�E���d�A}��������R�2��v�X,��>�ϊ}-C	$�V�	,1�L�"�@�
��BC��ep
Z��ڧV	�I�Dw�Ĺ| ��\�'i8��m�p��S�W�^�O����cV�(���:�GR:o��kޚ%'���E�ÄM�m�i�c¢���Y�M��'F�F�K>n"�c�,p�Ԥo�)5�m�P�+�֝��Bt�:�UO���g:�CV!�2�p���'9m��8D($]P�b�V@j2R�0wD��2��R��QP�SDJh�`!
���+
h_ `D�B3���+V�H�Qt��Ip&�q��x�/2p���I�X�|�2l�K%�|��d��2���䊕���$�*��v�T��<'x�7�,�d3E��/](\�����p���x�t~��,���������i�3�V���si��Ԗu�)��������Z�uBt�.h��Tɶѵ4I�{rǻCE*C��m�eD�=tn�Ʊ:�&�Q��w$S�	ռE�